----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:34:26 10/07/2016 
-- Design Name: 
-- Module Name:    nextProgramCounter - arq_nextProgramCounter 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use IEEE.STD_LOGIC_arith.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity nextProgramCounter is
    Port ( InAddress : in  STD_LOGIC_VECTOR (31 downto 0);
           clk : in  STD_LOGIC;
           Reset : in  STD_LOGIC;
           outAddress : out  STD_LOGIC_VECTOR (31 downto 0));
end nextProgramCounter;

architecture arq_nextProgramCounter of nextProgramCounter is

begin
	process(clk,Reset)

	begin

		if Reset = '1' then 
			OutAddress <= "00000000000000000000000000000000";
		elsif rising_edge(clk) then 
			OutAddress <= InAddress;
		end if;
	end process;

end arq_nextProgramCounter;

